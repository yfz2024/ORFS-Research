VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_2048x39_bottom
  FOREIGN fakeram45_2048x39_bottom 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 206.910 BY 219.800 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.800 0.070 2.870 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.200 0.070 4.270 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.600 0.070 5.670 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.000 0.070 7.070 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.400 0.070 8.470 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.800 0.070 9.870 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.200 0.070 11.270 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.600 0.070 12.670 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.000 0.070 14.070 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.400 0.070 15.470 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.800 0.070 16.870 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.200 0.070 18.270 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.600 0.070 19.670 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.000 0.070 21.070 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.400 0.070 22.470 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.800 0.070 23.870 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.200 0.070 25.270 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.600 0.070 26.670 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.000 0.070 28.070 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.400 0.070 29.470 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.800 0.070 30.870 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.200 0.070 32.270 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.600 0.070 33.670 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.000 0.070 35.070 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.400 0.070 36.470 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.800 0.070 37.870 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.200 0.070 39.270 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.600 0.070 40.670 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.000 0.070 42.070 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.400 0.070 43.470 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.800 0.070 44.870 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.200 0.070 46.270 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.600 0.070 47.670 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.000 0.070 49.070 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.400 0.070 50.470 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.800 0.070 51.870 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.200 0.070 53.270 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.600 0.070 54.670 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.000 0.070 56.070 ;
    END
  END w_mask_in[38]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.560 0.070 63.630 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.960 0.070 65.030 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.360 0.070 66.430 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.760 0.070 67.830 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.160 0.070 69.230 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.560 0.070 70.630 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.960 0.070 72.030 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.360 0.070 73.430 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.760 0.070 74.830 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.160 0.070 76.230 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.560 0.070 77.630 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.960 0.070 79.030 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.360 0.070 80.430 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.760 0.070 81.830 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.160 0.070 83.230 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.560 0.070 84.630 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.960 0.070 86.030 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.360 0.070 87.430 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.760 0.070 88.830 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.160 0.070 90.230 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.560 0.070 91.630 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.960 0.070 93.030 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.360 0.070 94.430 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.760 0.070 95.830 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.160 0.070 97.230 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.560 0.070 98.630 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.960 0.070 100.030 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.360 0.070 101.430 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.760 0.070 102.830 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.160 0.070 104.230 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.560 0.070 105.630 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.960 0.070 107.030 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.360 0.070 108.430 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.760 0.070 109.830 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.160 0.070 111.230 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.560 0.070 112.630 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.960 0.070 114.030 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.360 0.070 115.430 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.760 0.070 116.830 ;
    END
  END rd_out[38]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.320 0.070 124.390 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.720 0.070 125.790 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.120 0.070 127.190 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.520 0.070 128.590 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.920 0.070 129.990 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.320 0.070 131.390 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.720 0.070 132.790 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.120 0.070 134.190 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.520 0.070 135.590 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.920 0.070 136.990 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.320 0.070 138.390 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.720 0.070 139.790 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.120 0.070 141.190 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.520 0.070 142.590 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.920 0.070 143.990 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.320 0.070 145.390 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.720 0.070 146.790 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.120 0.070 148.190 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.520 0.070 149.590 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.920 0.070 150.990 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.320 0.070 152.390 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.720 0.070 153.790 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.120 0.070 155.190 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.520 0.070 156.590 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.920 0.070 157.990 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.320 0.070 159.390 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.720 0.070 160.790 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.120 0.070 162.190 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.520 0.070 163.590 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.920 0.070 164.990 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.320 0.070 166.390 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.720 0.070 167.790 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.120 0.070 169.190 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.520 0.070 170.590 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.920 0.070 171.990 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.320 0.070 173.390 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.720 0.070 174.790 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.120 0.070 176.190 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.520 0.070 177.590 ;
    END
  END wd_in[38]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.080 0.070 185.150 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.480 0.070 186.550 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.880 0.070 187.950 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.280 0.070 189.350 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.680 0.070 190.750 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.080 0.070 192.150 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.480 0.070 193.550 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.880 0.070 194.950 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.280 0.070 196.350 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.680 0.070 197.750 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.080 0.070 199.150 ;
    END
  END addr_in[10]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.640 0.070 206.710 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.040 0.070 208.110 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.440 0.070 209.510 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 2.660 2.800 2.940 217.000 ;
      RECT 7.140 2.800 7.420 217.000 ;
      RECT 11.620 2.800 11.900 217.000 ;
      RECT 16.100 2.800 16.380 217.000 ;
      RECT 20.580 2.800 20.860 217.000 ;
      RECT 25.060 2.800 25.340 217.000 ;
      RECT 29.540 2.800 29.820 217.000 ;
      RECT 34.020 2.800 34.300 217.000 ;
      RECT 38.500 2.800 38.780 217.000 ;
      RECT 42.980 2.800 43.260 217.000 ;
      RECT 47.460 2.800 47.740 217.000 ;
      RECT 51.940 2.800 52.220 217.000 ;
      RECT 56.420 2.800 56.700 217.000 ;
      RECT 60.900 2.800 61.180 217.000 ;
      RECT 65.380 2.800 65.660 217.000 ;
      RECT 69.860 2.800 70.140 217.000 ;
      RECT 74.340 2.800 74.620 217.000 ;
      RECT 78.820 2.800 79.100 217.000 ;
      RECT 83.300 2.800 83.580 217.000 ;
      RECT 87.780 2.800 88.060 217.000 ;
      RECT 92.260 2.800 92.540 217.000 ;
      RECT 96.740 2.800 97.020 217.000 ;
      RECT 101.220 2.800 101.500 217.000 ;
      RECT 105.700 2.800 105.980 217.000 ;
      RECT 110.180 2.800 110.460 217.000 ;
      RECT 114.660 2.800 114.940 217.000 ;
      RECT 119.140 2.800 119.420 217.000 ;
      RECT 123.620 2.800 123.900 217.000 ;
      RECT 128.100 2.800 128.380 217.000 ;
      RECT 132.580 2.800 132.860 217.000 ;
      RECT 137.060 2.800 137.340 217.000 ;
      RECT 141.540 2.800 141.820 217.000 ;
      RECT 146.020 2.800 146.300 217.000 ;
      RECT 150.500 2.800 150.780 217.000 ;
      RECT 154.980 2.800 155.260 217.000 ;
      RECT 159.460 2.800 159.740 217.000 ;
      RECT 163.940 2.800 164.220 217.000 ;
      RECT 168.420 2.800 168.700 217.000 ;
      RECT 172.900 2.800 173.180 217.000 ;
      RECT 177.380 2.800 177.660 217.000 ;
      RECT 181.860 2.800 182.140 217.000 ;
      RECT 186.340 2.800 186.620 217.000 ;
      RECT 190.820 2.800 191.100 217.000 ;
      RECT 195.300 2.800 195.580 217.000 ;
      RECT 199.780 2.800 200.060 217.000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 4.900 2.800 5.180 217.000 ;
      RECT 9.380 2.800 9.660 217.000 ;
      RECT 13.860 2.800 14.140 217.000 ;
      RECT 18.340 2.800 18.620 217.000 ;
      RECT 22.820 2.800 23.100 217.000 ;
      RECT 27.300 2.800 27.580 217.000 ;
      RECT 31.780 2.800 32.060 217.000 ;
      RECT 36.260 2.800 36.540 217.000 ;
      RECT 40.740 2.800 41.020 217.000 ;
      RECT 45.220 2.800 45.500 217.000 ;
      RECT 49.700 2.800 49.980 217.000 ;
      RECT 54.180 2.800 54.460 217.000 ;
      RECT 58.660 2.800 58.940 217.000 ;
      RECT 63.140 2.800 63.420 217.000 ;
      RECT 67.620 2.800 67.900 217.000 ;
      RECT 72.100 2.800 72.380 217.000 ;
      RECT 76.580 2.800 76.860 217.000 ;
      RECT 81.060 2.800 81.340 217.000 ;
      RECT 85.540 2.800 85.820 217.000 ;
      RECT 90.020 2.800 90.300 217.000 ;
      RECT 94.500 2.800 94.780 217.000 ;
      RECT 98.980 2.800 99.260 217.000 ;
      RECT 103.460 2.800 103.740 217.000 ;
      RECT 107.940 2.800 108.220 217.000 ;
      RECT 112.420 2.800 112.700 217.000 ;
      RECT 116.900 2.800 117.180 217.000 ;
      RECT 121.380 2.800 121.660 217.000 ;
      RECT 125.860 2.800 126.140 217.000 ;
      RECT 130.340 2.800 130.620 217.000 ;
      RECT 134.820 2.800 135.100 217.000 ;
      RECT 139.300 2.800 139.580 217.000 ;
      RECT 143.780 2.800 144.060 217.000 ;
      RECT 148.260 2.800 148.540 217.000 ;
      RECT 152.740 2.800 153.020 217.000 ;
      RECT 157.220 2.800 157.500 217.000 ;
      RECT 161.700 2.800 161.980 217.000 ;
      RECT 166.180 2.800 166.460 217.000 ;
      RECT 170.660 2.800 170.940 217.000 ;
      RECT 175.140 2.800 175.420 217.000 ;
      RECT 179.620 2.800 179.900 217.000 ;
      RECT 184.100 2.800 184.380 217.000 ;
      RECT 188.580 2.800 188.860 217.000 ;
      RECT 193.060 2.800 193.340 217.000 ;
      RECT 197.540 2.800 197.820 217.000 ;
      RECT 202.020 2.800 202.300 217.000 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 206.910 219.800 ;
    LAYER metal2 ;
    RECT 0 0 206.910 219.800 ;
    LAYER metal3 ;
    RECT 0.070 0 206.910 219.800 ;
    RECT 0 0.000 0.070 2.800 ;
    RECT 0 2.870 0.070 4.200 ;
    RECT 0 4.270 0.070 5.600 ;
    RECT 0 5.670 0.070 7.000 ;
    RECT 0 7.070 0.070 8.400 ;
    RECT 0 8.470 0.070 9.800 ;
    RECT 0 9.870 0.070 11.200 ;
    RECT 0 11.270 0.070 12.600 ;
    RECT 0 12.670 0.070 14.000 ;
    RECT 0 14.070 0.070 15.400 ;
    RECT 0 15.470 0.070 16.800 ;
    RECT 0 16.870 0.070 18.200 ;
    RECT 0 18.270 0.070 19.600 ;
    RECT 0 19.670 0.070 21.000 ;
    RECT 0 21.070 0.070 22.400 ;
    RECT 0 22.470 0.070 23.800 ;
    RECT 0 23.870 0.070 25.200 ;
    RECT 0 25.270 0.070 26.600 ;
    RECT 0 26.670 0.070 28.000 ;
    RECT 0 28.070 0.070 29.400 ;
    RECT 0 29.470 0.070 30.800 ;
    RECT 0 30.870 0.070 32.200 ;
    RECT 0 32.270 0.070 33.600 ;
    RECT 0 33.670 0.070 35.000 ;
    RECT 0 35.070 0.070 36.400 ;
    RECT 0 36.470 0.070 37.800 ;
    RECT 0 37.870 0.070 39.200 ;
    RECT 0 39.270 0.070 40.600 ;
    RECT 0 40.670 0.070 42.000 ;
    RECT 0 42.070 0.070 43.400 ;
    RECT 0 43.470 0.070 44.800 ;
    RECT 0 44.870 0.070 46.200 ;
    RECT 0 46.270 0.070 47.600 ;
    RECT 0 47.670 0.070 49.000 ;
    RECT 0 49.070 0.070 50.400 ;
    RECT 0 50.470 0.070 51.800 ;
    RECT 0 51.870 0.070 53.200 ;
    RECT 0 53.270 0.070 54.600 ;
    RECT 0 54.670 0.070 56.000 ;
    RECT 0 56.070 0.070 63.560 ;
    RECT 0 63.630 0.070 64.960 ;
    RECT 0 65.030 0.070 66.360 ;
    RECT 0 66.430 0.070 67.760 ;
    RECT 0 67.830 0.070 69.160 ;
    RECT 0 69.230 0.070 70.560 ;
    RECT 0 70.630 0.070 71.960 ;
    RECT 0 72.030 0.070 73.360 ;
    RECT 0 73.430 0.070 74.760 ;
    RECT 0 74.830 0.070 76.160 ;
    RECT 0 76.230 0.070 77.560 ;
    RECT 0 77.630 0.070 78.960 ;
    RECT 0 79.030 0.070 80.360 ;
    RECT 0 80.430 0.070 81.760 ;
    RECT 0 81.830 0.070 83.160 ;
    RECT 0 83.230 0.070 84.560 ;
    RECT 0 84.630 0.070 85.960 ;
    RECT 0 86.030 0.070 87.360 ;
    RECT 0 87.430 0.070 88.760 ;
    RECT 0 88.830 0.070 90.160 ;
    RECT 0 90.230 0.070 91.560 ;
    RECT 0 91.630 0.070 92.960 ;
    RECT 0 93.030 0.070 94.360 ;
    RECT 0 94.430 0.070 95.760 ;
    RECT 0 95.830 0.070 97.160 ;
    RECT 0 97.230 0.070 98.560 ;
    RECT 0 98.630 0.070 99.960 ;
    RECT 0 100.030 0.070 101.360 ;
    RECT 0 101.430 0.070 102.760 ;
    RECT 0 102.830 0.070 104.160 ;
    RECT 0 104.230 0.070 105.560 ;
    RECT 0 105.630 0.070 106.960 ;
    RECT 0 107.030 0.070 108.360 ;
    RECT 0 108.430 0.070 109.760 ;
    RECT 0 109.830 0.070 111.160 ;
    RECT 0 111.230 0.070 112.560 ;
    RECT 0 112.630 0.070 113.960 ;
    RECT 0 114.030 0.070 115.360 ;
    RECT 0 115.430 0.070 116.760 ;
    RECT 0 116.830 0.070 124.320 ;
    RECT 0 124.390 0.070 125.720 ;
    RECT 0 125.790 0.070 127.120 ;
    RECT 0 127.190 0.070 128.520 ;
    RECT 0 128.590 0.070 129.920 ;
    RECT 0 129.990 0.070 131.320 ;
    RECT 0 131.390 0.070 132.720 ;
    RECT 0 132.790 0.070 134.120 ;
    RECT 0 134.190 0.070 135.520 ;
    RECT 0 135.590 0.070 136.920 ;
    RECT 0 136.990 0.070 138.320 ;
    RECT 0 138.390 0.070 139.720 ;
    RECT 0 139.790 0.070 141.120 ;
    RECT 0 141.190 0.070 142.520 ;
    RECT 0 142.590 0.070 143.920 ;
    RECT 0 143.990 0.070 145.320 ;
    RECT 0 145.390 0.070 146.720 ;
    RECT 0 146.790 0.070 148.120 ;
    RECT 0 148.190 0.070 149.520 ;
    RECT 0 149.590 0.070 150.920 ;
    RECT 0 150.990 0.070 152.320 ;
    RECT 0 152.390 0.070 153.720 ;
    RECT 0 153.790 0.070 155.120 ;
    RECT 0 155.190 0.070 156.520 ;
    RECT 0 156.590 0.070 157.920 ;
    RECT 0 157.990 0.070 159.320 ;
    RECT 0 159.390 0.070 160.720 ;
    RECT 0 160.790 0.070 162.120 ;
    RECT 0 162.190 0.070 163.520 ;
    RECT 0 163.590 0.070 164.920 ;
    RECT 0 164.990 0.070 166.320 ;
    RECT 0 166.390 0.070 167.720 ;
    RECT 0 167.790 0.070 169.120 ;
    RECT 0 169.190 0.070 170.520 ;
    RECT 0 170.590 0.070 171.920 ;
    RECT 0 171.990 0.070 173.320 ;
    RECT 0 173.390 0.070 174.720 ;
    RECT 0 174.790 0.070 176.120 ;
    RECT 0 176.190 0.070 177.520 ;
    RECT 0 177.590 0.070 185.080 ;
    RECT 0 185.150 0.070 186.480 ;
    RECT 0 186.550 0.070 187.880 ;
    RECT 0 187.950 0.070 189.280 ;
    RECT 0 189.350 0.070 190.680 ;
    RECT 0 190.750 0.070 192.080 ;
    RECT 0 192.150 0.070 193.480 ;
    RECT 0 193.550 0.070 194.880 ;
    RECT 0 194.950 0.070 196.280 ;
    RECT 0 196.350 0.070 197.680 ;
    RECT 0 197.750 0.070 199.080 ;
    RECT 0 199.150 0.070 206.640 ;
    RECT 0 206.710 0.070 208.040 ;
    RECT 0 208.110 0.070 209.440 ;
    RECT 0 209.510 0.070 219.800 ;
    LAYER metal4 ;
    RECT 0 0 206.910 2.800 ;
    RECT 0 217.000 206.910 219.800 ;
    RECT 0.000 2.800 2.660 217.000 ;
    RECT 2.940 2.800 4.900 217.000 ;
    RECT 5.180 2.800 7.140 217.000 ;
    RECT 7.420 2.800 9.380 217.000 ;
    RECT 9.660 2.800 11.620 217.000 ;
    RECT 11.900 2.800 13.860 217.000 ;
    RECT 14.140 2.800 16.100 217.000 ;
    RECT 16.380 2.800 18.340 217.000 ;
    RECT 18.620 2.800 20.580 217.000 ;
    RECT 20.860 2.800 22.820 217.000 ;
    RECT 23.100 2.800 25.060 217.000 ;
    RECT 25.340 2.800 27.300 217.000 ;
    RECT 27.580 2.800 29.540 217.000 ;
    RECT 29.820 2.800 31.780 217.000 ;
    RECT 32.060 2.800 34.020 217.000 ;
    RECT 34.300 2.800 36.260 217.000 ;
    RECT 36.540 2.800 38.500 217.000 ;
    RECT 38.780 2.800 40.740 217.000 ;
    RECT 41.020 2.800 42.980 217.000 ;
    RECT 43.260 2.800 45.220 217.000 ;
    RECT 45.500 2.800 47.460 217.000 ;
    RECT 47.740 2.800 49.700 217.000 ;
    RECT 49.980 2.800 51.940 217.000 ;
    RECT 52.220 2.800 54.180 217.000 ;
    RECT 54.460 2.800 56.420 217.000 ;
    RECT 56.700 2.800 58.660 217.000 ;
    RECT 58.940 2.800 60.900 217.000 ;
    RECT 61.180 2.800 63.140 217.000 ;
    RECT 63.420 2.800 65.380 217.000 ;
    RECT 65.660 2.800 67.620 217.000 ;
    RECT 67.900 2.800 69.860 217.000 ;
    RECT 70.140 2.800 72.100 217.000 ;
    RECT 72.380 2.800 74.340 217.000 ;
    RECT 74.620 2.800 76.580 217.000 ;
    RECT 76.860 2.800 78.820 217.000 ;
    RECT 79.100 2.800 81.060 217.000 ;
    RECT 81.340 2.800 83.300 217.000 ;
    RECT 83.580 2.800 85.540 217.000 ;
    RECT 85.820 2.800 87.780 217.000 ;
    RECT 88.060 2.800 90.020 217.000 ;
    RECT 90.300 2.800 92.260 217.000 ;
    RECT 92.540 2.800 94.500 217.000 ;
    RECT 94.780 2.800 96.740 217.000 ;
    RECT 97.020 2.800 98.980 217.000 ;
    RECT 99.260 2.800 101.220 217.000 ;
    RECT 101.500 2.800 103.460 217.000 ;
    RECT 103.740 2.800 105.700 217.000 ;
    RECT 105.980 2.800 107.940 217.000 ;
    RECT 108.220 2.800 110.180 217.000 ;
    RECT 110.460 2.800 112.420 217.000 ;
    RECT 112.700 2.800 114.660 217.000 ;
    RECT 114.940 2.800 116.900 217.000 ;
    RECT 117.180 2.800 119.140 217.000 ;
    RECT 119.420 2.800 121.380 217.000 ;
    RECT 121.660 2.800 123.620 217.000 ;
    RECT 123.900 2.800 125.860 217.000 ;
    RECT 126.140 2.800 128.100 217.000 ;
    RECT 128.380 2.800 130.340 217.000 ;
    RECT 130.620 2.800 132.580 217.000 ;
    RECT 132.860 2.800 134.820 217.000 ;
    RECT 135.100 2.800 137.060 217.000 ;
    RECT 137.340 2.800 139.300 217.000 ;
    RECT 139.580 2.800 141.540 217.000 ;
    RECT 141.820 2.800 143.780 217.000 ;
    RECT 144.060 2.800 146.020 217.000 ;
    RECT 146.300 2.800 148.260 217.000 ;
    RECT 148.540 2.800 150.500 217.000 ;
    RECT 150.780 2.800 152.740 217.000 ;
    RECT 153.020 2.800 154.980 217.000 ;
    RECT 155.260 2.800 157.220 217.000 ;
    RECT 157.500 2.800 159.460 217.000 ;
    RECT 159.740 2.800 161.700 217.000 ;
    RECT 161.980 2.800 163.940 217.000 ;
    RECT 164.220 2.800 166.180 217.000 ;
    RECT 166.460 2.800 168.420 217.000 ;
    RECT 168.700 2.800 170.660 217.000 ;
    RECT 170.940 2.800 172.900 217.000 ;
    RECT 173.180 2.800 175.140 217.000 ;
    RECT 175.420 2.800 177.380 217.000 ;
    RECT 177.660 2.800 179.620 217.000 ;
    RECT 179.900 2.800 181.860 217.000 ;
    RECT 182.140 2.800 184.100 217.000 ;
    RECT 184.380 2.800 186.340 217.000 ;
    RECT 186.620 2.800 188.580 217.000 ;
    RECT 188.860 2.800 190.820 217.000 ;
    RECT 191.100 2.800 193.060 217.000 ;
    RECT 193.340 2.800 195.300 217.000 ;
    RECT 195.580 2.800 197.540 217.000 ;
    RECT 197.820 2.800 199.780 217.000 ;
    RECT 200.060 2.800 202.020 217.000 ;
    RECT 202.300 2.800 206.910 217.000 ;
  END
END fakeram45_2048x39_bottom

END LIBRARY
