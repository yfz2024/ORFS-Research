VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_64x64_upper
  FOREIGN fakeram45_64x64_upper 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 77.900 BY 62.200 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 2.800 0.070 2.870 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 3.080 0.070 3.150 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 3.360 0.070 3.430 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 3.640 0.070 3.710 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 3.920 0.070 3.990 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 4.200 0.070 4.270 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 4.480 0.070 4.550 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 4.760 0.070 4.830 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 5.040 0.070 5.110 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 5.320 0.070 5.390 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 5.600 0.070 5.670 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 5.880 0.070 5.950 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 6.160 0.070 6.230 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 6.440 0.070 6.510 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 6.720 0.070 6.790 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 7.000 0.070 7.070 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 7.280 0.070 7.350 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 7.560 0.070 7.630 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 7.840 0.070 7.910 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 8.120 0.070 8.190 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 8.400 0.070 8.470 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 8.680 0.070 8.750 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 8.960 0.070 9.030 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 9.240 0.070 9.310 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 9.520 0.070 9.590 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 9.800 0.070 9.870 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 10.080 0.070 10.150 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 10.360 0.070 10.430 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 10.640 0.070 10.710 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 10.920 0.070 10.990 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 11.200 0.070 11.270 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 11.480 0.070 11.550 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 11.760 0.070 11.830 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 12.040 0.070 12.110 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 12.320 0.070 12.390 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 12.600 0.070 12.670 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 12.880 0.070 12.950 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 13.160 0.070 13.230 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 13.440 0.070 13.510 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 13.720 0.070 13.790 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 14.000 0.070 14.070 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 14.280 0.070 14.350 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 14.560 0.070 14.630 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 14.840 0.070 14.910 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 15.120 0.070 15.190 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 15.400 0.070 15.470 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 15.680 0.070 15.750 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 15.960 0.070 16.030 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 16.240 0.070 16.310 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 16.520 0.070 16.590 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 16.800 0.070 16.870 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 17.080 0.070 17.150 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 17.360 0.070 17.430 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 17.640 0.070 17.710 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 17.920 0.070 17.990 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 18.200 0.070 18.270 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 18.480 0.070 18.550 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 18.760 0.070 18.830 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 19.040 0.070 19.110 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 19.320 0.070 19.390 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 19.600 0.070 19.670 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 19.880 0.070 19.950 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 20.160 0.070 20.230 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 20.440 0.070 20.510 ;
    END
  END w_mask_in[63]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 20.720 0.070 20.790 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 21.000 0.070 21.070 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 21.280 0.070 21.350 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 21.560 0.070 21.630 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 21.840 0.070 21.910 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 22.120 0.070 22.190 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 22.400 0.070 22.470 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 22.680 0.070 22.750 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 22.960 0.070 23.030 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 23.240 0.070 23.310 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 23.520 0.070 23.590 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 23.800 0.070 23.870 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 24.080 0.070 24.150 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 24.360 0.070 24.430 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 24.640 0.070 24.710 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 24.920 0.070 24.990 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 25.200 0.070 25.270 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 25.480 0.070 25.550 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 25.760 0.070 25.830 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 26.040 0.070 26.110 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 26.320 0.070 26.390 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 26.600 0.070 26.670 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 26.880 0.070 26.950 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 27.160 0.070 27.230 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 27.440 0.070 27.510 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 27.720 0.070 27.790 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 28.000 0.070 28.070 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 28.280 0.070 28.350 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 28.560 0.070 28.630 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 28.840 0.070 28.910 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 29.120 0.070 29.190 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 29.400 0.070 29.470 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 29.680 0.070 29.750 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 29.960 0.070 30.030 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 30.240 0.070 30.310 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 30.520 0.070 30.590 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 30.800 0.070 30.870 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 31.080 0.070 31.150 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 31.360 0.070 31.430 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 31.640 0.070 31.710 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 31.920 0.070 31.990 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 32.200 0.070 32.270 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 32.480 0.070 32.550 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 32.760 0.070 32.830 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 33.040 0.070 33.110 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 33.320 0.070 33.390 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 33.600 0.070 33.670 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 33.880 0.070 33.950 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 34.160 0.070 34.230 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 34.440 0.070 34.510 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 34.720 0.070 34.790 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 35.000 0.070 35.070 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 35.280 0.070 35.350 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 35.560 0.070 35.630 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 35.840 0.070 35.910 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 36.120 0.070 36.190 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 36.400 0.070 36.470 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 36.680 0.070 36.750 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 36.960 0.070 37.030 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 37.240 0.070 37.310 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 37.520 0.070 37.590 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 37.800 0.070 37.870 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 38.080 0.070 38.150 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 38.360 0.070 38.430 ;
    END
  END rd_out[63]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 38.640 0.070 38.710 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 38.920 0.070 38.990 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 39.200 0.070 39.270 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 39.480 0.070 39.550 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 39.760 0.070 39.830 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 40.040 0.070 40.110 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 40.320 0.070 40.390 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 40.600 0.070 40.670 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 40.880 0.070 40.950 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 41.160 0.070 41.230 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 41.440 0.070 41.510 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 41.720 0.070 41.790 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 42.000 0.070 42.070 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 42.280 0.070 42.350 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 42.560 0.070 42.630 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 42.840 0.070 42.910 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 43.120 0.070 43.190 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 43.400 0.070 43.470 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 43.680 0.070 43.750 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 43.960 0.070 44.030 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 44.240 0.070 44.310 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 44.520 0.070 44.590 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 44.800 0.070 44.870 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 45.080 0.070 45.150 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 45.360 0.070 45.430 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 45.640 0.070 45.710 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 45.920 0.070 45.990 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 46.200 0.070 46.270 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 46.480 0.070 46.550 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 46.760 0.070 46.830 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 47.040 0.070 47.110 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 47.320 0.070 47.390 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 47.600 0.070 47.670 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 47.880 0.070 47.950 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 48.160 0.070 48.230 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 48.440 0.070 48.510 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 48.720 0.070 48.790 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 49.000 0.070 49.070 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 49.280 0.070 49.350 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 49.560 0.070 49.630 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 49.840 0.070 49.910 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 50.120 0.070 50.190 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 50.400 0.070 50.470 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 50.680 0.070 50.750 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 50.960 0.070 51.030 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 51.240 0.070 51.310 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 51.520 0.070 51.590 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 51.800 0.070 51.870 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 52.080 0.070 52.150 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 52.360 0.070 52.430 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 52.640 0.070 52.710 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 52.920 0.070 52.990 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 53.200 0.070 53.270 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 53.480 0.070 53.550 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 53.760 0.070 53.830 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 54.040 0.070 54.110 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 54.320 0.070 54.390 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 54.600 0.070 54.670 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 54.880 0.070 54.950 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 55.160 0.070 55.230 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 55.440 0.070 55.510 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 55.720 0.070 55.790 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 56.000 0.070 56.070 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 56.280 0.070 56.350 ;
    END
  END wd_in[63]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 56.560 0.070 56.630 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 56.840 0.070 56.910 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 57.120 0.070 57.190 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 57.400 0.070 57.470 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 57.680 0.070 57.750 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 57.960 0.070 58.030 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 58.240 0.070 58.310 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 58.520 0.070 58.590 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 58.800 0.070 58.870 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal17 ;
      RECT 2.660 2.800 2.940 59.400 ;
      RECT 7.140 2.800 7.420 59.400 ;
      RECT 11.620 2.800 11.900 59.400 ;
      RECT 16.100 2.800 16.380 59.400 ;
      RECT 20.580 2.800 20.860 59.400 ;
      RECT 25.060 2.800 25.340 59.400 ;
      RECT 29.540 2.800 29.820 59.400 ;
      RECT 34.020 2.800 34.300 59.400 ;
      RECT 38.500 2.800 38.780 59.400 ;
      RECT 42.980 2.800 43.260 59.400 ;
      RECT 47.460 2.800 47.740 59.400 ;
      RECT 51.940 2.800 52.220 59.400 ;
      RECT 56.420 2.800 56.700 59.400 ;
      RECT 60.900 2.800 61.180 59.400 ;
      RECT 65.380 2.800 65.660 59.400 ;
      RECT 69.860 2.800 70.140 59.400 ;
      RECT 74.340 2.800 74.620 59.400 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal17 ;
      RECT 4.900 2.800 5.180 59.400 ;
      RECT 9.380 2.800 9.660 59.400 ;
      RECT 13.860 2.800 14.140 59.400 ;
      RECT 18.340 2.800 18.620 59.400 ;
      RECT 22.820 2.800 23.100 59.400 ;
      RECT 27.300 2.800 27.580 59.400 ;
      RECT 31.780 2.800 32.060 59.400 ;
      RECT 36.260 2.800 36.540 59.400 ;
      RECT 40.740 2.800 41.020 59.400 ;
      RECT 45.220 2.800 45.500 59.400 ;
      RECT 49.700 2.800 49.980 59.400 ;
      RECT 54.180 2.800 54.460 59.400 ;
      RECT 58.660 2.800 58.940 59.400 ;
      RECT 63.140 2.800 63.420 59.400 ;
      RECT 67.620 2.800 67.900 59.400 ;
      RECT 72.100 2.800 72.380 59.400 ;
    END
  END VDD
  OBS
    LAYER metal20 ;
    RECT 0 0 77.900 62.200 ;
    LAYER metal19 ;
    RECT 0 0 77.900 62.200 ;
    LAYER metal18 ;
    RECT 0.070 0 77.900 62.200 ;
    RECT 0 0.000 0.070 2.800 ;
    RECT 0 2.870 0.070 3.080 ;
    RECT 0 3.150 0.070 3.360 ;
    RECT 0 3.430 0.070 3.640 ;
    RECT 0 3.710 0.070 3.920 ;
    RECT 0 3.990 0.070 4.200 ;
    RECT 0 4.270 0.070 4.480 ;
    RECT 0 4.550 0.070 4.760 ;
    RECT 0 4.830 0.070 5.040 ;
    RECT 0 5.110 0.070 5.320 ;
    RECT 0 5.390 0.070 5.600 ;
    RECT 0 5.670 0.070 5.880 ;
    RECT 0 5.950 0.070 6.160 ;
    RECT 0 6.230 0.070 6.440 ;
    RECT 0 6.510 0.070 6.720 ;
    RECT 0 6.790 0.070 7.000 ;
    RECT 0 7.070 0.070 7.280 ;
    RECT 0 7.350 0.070 7.560 ;
    RECT 0 7.630 0.070 7.840 ;
    RECT 0 7.910 0.070 8.120 ;
    RECT 0 8.190 0.070 8.400 ;
    RECT 0 8.470 0.070 8.680 ;
    RECT 0 8.750 0.070 8.960 ;
    RECT 0 9.030 0.070 9.240 ;
    RECT 0 9.310 0.070 9.520 ;
    RECT 0 9.590 0.070 9.800 ;
    RECT 0 9.870 0.070 10.080 ;
    RECT 0 10.150 0.070 10.360 ;
    RECT 0 10.430 0.070 10.640 ;
    RECT 0 10.710 0.070 10.920 ;
    RECT 0 10.990 0.070 11.200 ;
    RECT 0 11.270 0.070 11.480 ;
    RECT 0 11.550 0.070 11.760 ;
    RECT 0 11.830 0.070 12.040 ;
    RECT 0 12.110 0.070 12.320 ;
    RECT 0 12.390 0.070 12.600 ;
    RECT 0 12.670 0.070 12.880 ;
    RECT 0 12.950 0.070 13.160 ;
    RECT 0 13.230 0.070 13.440 ;
    RECT 0 13.510 0.070 13.720 ;
    RECT 0 13.790 0.070 14.000 ;
    RECT 0 14.070 0.070 14.280 ;
    RECT 0 14.350 0.070 14.560 ;
    RECT 0 14.630 0.070 14.840 ;
    RECT 0 14.910 0.070 15.120 ;
    RECT 0 15.190 0.070 15.400 ;
    RECT 0 15.470 0.070 15.680 ;
    RECT 0 15.750 0.070 15.960 ;
    RECT 0 16.030 0.070 16.240 ;
    RECT 0 16.310 0.070 16.520 ;
    RECT 0 16.590 0.070 16.800 ;
    RECT 0 16.870 0.070 17.080 ;
    RECT 0 17.150 0.070 17.360 ;
    RECT 0 17.430 0.070 17.640 ;
    RECT 0 17.710 0.070 17.920 ;
    RECT 0 17.990 0.070 18.200 ;
    RECT 0 18.270 0.070 18.480 ;
    RECT 0 18.550 0.070 18.760 ;
    RECT 0 18.830 0.070 19.040 ;
    RECT 0 19.110 0.070 19.320 ;
    RECT 0 19.390 0.070 19.600 ;
    RECT 0 19.670 0.070 19.880 ;
    RECT 0 19.950 0.070 20.160 ;
    RECT 0 20.230 0.070 20.440 ;
    RECT 0 20.510 0.070 20.720 ;
    RECT 0 20.790 0.070 21.000 ;
    RECT 0 21.070 0.070 21.280 ;
    RECT 0 21.350 0.070 21.560 ;
    RECT 0 21.630 0.070 21.840 ;
    RECT 0 21.910 0.070 22.120 ;
    RECT 0 22.190 0.070 22.400 ;
    RECT 0 22.470 0.070 22.680 ;
    RECT 0 22.750 0.070 22.960 ;
    RECT 0 23.030 0.070 23.240 ;
    RECT 0 23.310 0.070 23.520 ;
    RECT 0 23.590 0.070 23.800 ;
    RECT 0 23.870 0.070 24.080 ;
    RECT 0 24.150 0.070 24.360 ;
    RECT 0 24.430 0.070 24.640 ;
    RECT 0 24.710 0.070 24.920 ;
    RECT 0 24.990 0.070 25.200 ;
    RECT 0 25.270 0.070 25.480 ;
    RECT 0 25.550 0.070 25.760 ;
    RECT 0 25.830 0.070 26.040 ;
    RECT 0 26.110 0.070 26.320 ;
    RECT 0 26.390 0.070 26.600 ;
    RECT 0 26.670 0.070 26.880 ;
    RECT 0 26.950 0.070 27.160 ;
    RECT 0 27.230 0.070 27.440 ;
    RECT 0 27.510 0.070 27.720 ;
    RECT 0 27.790 0.070 28.000 ;
    RECT 0 28.070 0.070 28.280 ;
    RECT 0 28.350 0.070 28.560 ;
    RECT 0 28.630 0.070 28.840 ;
    RECT 0 28.910 0.070 29.120 ;
    RECT 0 29.190 0.070 29.400 ;
    RECT 0 29.470 0.070 29.680 ;
    RECT 0 29.750 0.070 29.960 ;
    RECT 0 30.030 0.070 30.240 ;
    RECT 0 30.310 0.070 30.520 ;
    RECT 0 30.590 0.070 30.800 ;
    RECT 0 30.870 0.070 31.080 ;
    RECT 0 31.150 0.070 31.360 ;
    RECT 0 31.430 0.070 31.640 ;
    RECT 0 31.710 0.070 31.920 ;
    RECT 0 31.990 0.070 32.200 ;
    RECT 0 32.270 0.070 32.480 ;
    RECT 0 32.550 0.070 32.760 ;
    RECT 0 32.830 0.070 33.040 ;
    RECT 0 33.110 0.070 33.320 ;
    RECT 0 33.390 0.070 33.600 ;
    RECT 0 33.670 0.070 33.880 ;
    RECT 0 33.950 0.070 34.160 ;
    RECT 0 34.230 0.070 34.440 ;
    RECT 0 34.510 0.070 34.720 ;
    RECT 0 34.790 0.070 35.000 ;
    RECT 0 35.070 0.070 35.280 ;
    RECT 0 35.350 0.070 35.560 ;
    RECT 0 35.630 0.070 35.840 ;
    RECT 0 35.910 0.070 36.120 ;
    RECT 0 36.190 0.070 36.400 ;
    RECT 0 36.470 0.070 36.680 ;
    RECT 0 36.750 0.070 36.960 ;
    RECT 0 37.030 0.070 37.240 ;
    RECT 0 37.310 0.070 37.520 ;
    RECT 0 37.590 0.070 37.800 ;
    RECT 0 37.870 0.070 38.080 ;
    RECT 0 38.150 0.070 38.360 ;
    RECT 0 38.430 0.070 38.640 ;
    RECT 0 38.710 0.070 38.920 ;
    RECT 0 38.990 0.070 39.200 ;
    RECT 0 39.270 0.070 39.480 ;
    RECT 0 39.550 0.070 39.760 ;
    RECT 0 39.830 0.070 40.040 ;
    RECT 0 40.110 0.070 40.320 ;
    RECT 0 40.390 0.070 40.600 ;
    RECT 0 40.670 0.070 40.880 ;
    RECT 0 40.950 0.070 41.160 ;
    RECT 0 41.230 0.070 41.440 ;
    RECT 0 41.510 0.070 41.720 ;
    RECT 0 41.790 0.070 42.000 ;
    RECT 0 42.070 0.070 42.280 ;
    RECT 0 42.350 0.070 42.560 ;
    RECT 0 42.630 0.070 42.840 ;
    RECT 0 42.910 0.070 43.120 ;
    RECT 0 43.190 0.070 43.400 ;
    RECT 0 43.470 0.070 43.680 ;
    RECT 0 43.750 0.070 43.960 ;
    RECT 0 44.030 0.070 44.240 ;
    RECT 0 44.310 0.070 44.520 ;
    RECT 0 44.590 0.070 44.800 ;
    RECT 0 44.870 0.070 45.080 ;
    RECT 0 45.150 0.070 45.360 ;
    RECT 0 45.430 0.070 45.640 ;
    RECT 0 45.710 0.070 45.920 ;
    RECT 0 45.990 0.070 46.200 ;
    RECT 0 46.270 0.070 46.480 ;
    RECT 0 46.550 0.070 46.760 ;
    RECT 0 46.830 0.070 47.040 ;
    RECT 0 47.110 0.070 47.320 ;
    RECT 0 47.390 0.070 47.600 ;
    RECT 0 47.670 0.070 47.880 ;
    RECT 0 47.950 0.070 48.160 ;
    RECT 0 48.230 0.070 48.440 ;
    RECT 0 48.510 0.070 48.720 ;
    RECT 0 48.790 0.070 49.000 ;
    RECT 0 49.070 0.070 49.280 ;
    RECT 0 49.350 0.070 49.560 ;
    RECT 0 49.630 0.070 49.840 ;
    RECT 0 49.910 0.070 50.120 ;
    RECT 0 50.190 0.070 50.400 ;
    RECT 0 50.470 0.070 50.680 ;
    RECT 0 50.750 0.070 50.960 ;
    RECT 0 51.030 0.070 51.240 ;
    RECT 0 51.310 0.070 51.520 ;
    RECT 0 51.590 0.070 51.800 ;
    RECT 0 51.870 0.070 52.080 ;
    RECT 0 52.150 0.070 52.360 ;
    RECT 0 52.430 0.070 52.640 ;
    RECT 0 52.710 0.070 52.920 ;
    RECT 0 52.990 0.070 53.200 ;
    RECT 0 53.270 0.070 53.480 ;
    RECT 0 53.550 0.070 53.760 ;
    RECT 0 53.830 0.070 54.040 ;
    RECT 0 54.110 0.070 54.320 ;
    RECT 0 54.390 0.070 54.600 ;
    RECT 0 54.670 0.070 54.880 ;
    RECT 0 54.950 0.070 55.160 ;
    RECT 0 55.230 0.070 55.440 ;
    RECT 0 55.510 0.070 55.720 ;
    RECT 0 55.790 0.070 56.000 ;
    RECT 0 56.070 0.070 56.280 ;
    RECT 0 56.350 0.070 56.560 ;
    RECT 0 56.630 0.070 56.840 ;
    RECT 0 56.910 0.070 57.120 ;
    RECT 0 57.190 0.070 57.400 ;
    RECT 0 57.470 0.070 57.680 ;
    RECT 0 57.750 0.070 57.960 ;
    RECT 0 58.030 0.070 58.240 ;
    RECT 0 58.310 0.070 58.520 ;
    RECT 0 58.590 0.070 58.800 ;
    RECT 0 58.870 0.070 62.200 ;
    LAYER metal17 ;
    RECT 0 0 77.900 2.800 ;
    RECT 0 59.400 77.900 62.200 ;
    RECT 0.000 2.800 2.660 59.400 ;
    RECT 2.940 2.800 4.900 59.400 ;
    RECT 5.180 2.800 7.140 59.400 ;
    RECT 7.420 2.800 9.380 59.400 ;
    RECT 9.660 2.800 11.620 59.400 ;
    RECT 11.900 2.800 13.860 59.400 ;
    RECT 14.140 2.800 16.100 59.400 ;
    RECT 16.380 2.800 18.340 59.400 ;
    RECT 18.620 2.800 20.580 59.400 ;
    RECT 20.860 2.800 22.820 59.400 ;
    RECT 23.100 2.800 25.060 59.400 ;
    RECT 25.340 2.800 27.300 59.400 ;
    RECT 27.580 2.800 29.540 59.400 ;
    RECT 29.820 2.800 31.780 59.400 ;
    RECT 32.060 2.800 34.020 59.400 ;
    RECT 34.300 2.800 36.260 59.400 ;
    RECT 36.540 2.800 38.500 59.400 ;
    RECT 38.780 2.800 40.740 59.400 ;
    RECT 41.020 2.800 42.980 59.400 ;
    RECT 43.260 2.800 45.220 59.400 ;
    RECT 45.500 2.800 47.460 59.400 ;
    RECT 47.740 2.800 49.700 59.400 ;
    RECT 49.980 2.800 51.940 59.400 ;
    RECT 52.220 2.800 54.180 59.400 ;
    RECT 54.460 2.800 56.420 59.400 ;
    RECT 56.700 2.800 58.660 59.400 ;
    RECT 58.940 2.800 60.900 59.400 ;
    RECT 61.180 2.800 63.140 59.400 ;
    RECT 63.420 2.800 65.380 59.400 ;
    RECT 65.660 2.800 67.620 59.400 ;
    RECT 67.900 2.800 69.860 59.400 ;
    RECT 70.140 2.800 72.100 59.400 ;
    RECT 72.380 2.800 74.340 59.400 ;
    RECT 74.620 2.800 77.900 59.400 ;
  END
END fakeram45_64x64_upper

END LIBRARY
