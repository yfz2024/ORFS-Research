VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_64x32_upper
  FOREIGN fakeram45_64x32_upper 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 20.140 BY 61.600 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 2.800 0.070 2.870 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 3.080 0.070 3.150 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 3.360 0.070 3.430 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 3.640 0.070 3.710 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 3.920 0.070 3.990 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 4.200 0.070 4.270 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 4.480 0.070 4.550 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 4.760 0.070 4.830 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 5.040 0.070 5.110 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 5.320 0.070 5.390 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 5.600 0.070 5.670 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 5.880 0.070 5.950 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 6.160 0.070 6.230 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 6.440 0.070 6.510 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 6.720 0.070 6.790 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 7.000 0.070 7.070 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 7.280 0.070 7.350 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 7.560 0.070 7.630 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 7.840 0.070 7.910 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 8.120 0.070 8.190 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 8.400 0.070 8.470 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 8.680 0.070 8.750 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 8.960 0.070 9.030 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 9.240 0.070 9.310 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 9.520 0.070 9.590 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 9.800 0.070 9.870 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 10.080 0.070 10.150 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 10.360 0.070 10.430 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 10.640 0.070 10.710 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 10.920 0.070 10.990 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 11.200 0.070 11.270 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 11.480 0.070 11.550 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 17.920 0.070 17.990 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 18.200 0.070 18.270 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 18.480 0.070 18.550 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 18.760 0.070 18.830 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 19.040 0.070 19.110 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 19.320 0.070 19.390 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 19.600 0.070 19.670 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 19.880 0.070 19.950 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 20.160 0.070 20.230 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 20.440 0.070 20.510 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 20.720 0.070 20.790 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 21.000 0.070 21.070 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 21.280 0.070 21.350 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 21.560 0.070 21.630 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 21.840 0.070 21.910 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 22.120 0.070 22.190 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 22.400 0.070 22.470 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 22.680 0.070 22.750 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 22.960 0.070 23.030 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 23.240 0.070 23.310 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 23.520 0.070 23.590 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 23.800 0.070 23.870 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 24.080 0.070 24.150 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 24.360 0.070 24.430 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 24.640 0.070 24.710 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 24.920 0.070 24.990 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 25.200 0.070 25.270 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 25.480 0.070 25.550 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 25.760 0.070 25.830 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 26.040 0.070 26.110 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 26.320 0.070 26.390 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 26.600 0.070 26.670 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 33.040 0.070 33.110 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 33.320 0.070 33.390 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 33.600 0.070 33.670 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 33.880 0.070 33.950 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 34.160 0.070 34.230 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 34.440 0.070 34.510 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 34.720 0.070 34.790 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 35.000 0.070 35.070 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 35.280 0.070 35.350 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 35.560 0.070 35.630 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 35.840 0.070 35.910 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 36.120 0.070 36.190 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 36.400 0.070 36.470 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 36.680 0.070 36.750 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 36.960 0.070 37.030 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 37.240 0.070 37.310 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 37.520 0.070 37.590 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 37.800 0.070 37.870 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 38.080 0.070 38.150 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 38.360 0.070 38.430 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 38.640 0.070 38.710 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 38.920 0.070 38.990 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 39.200 0.070 39.270 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 39.480 0.070 39.550 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 39.760 0.070 39.830 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 40.040 0.070 40.110 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 40.320 0.070 40.390 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 40.600 0.070 40.670 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 40.880 0.070 40.950 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 41.160 0.070 41.230 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 41.440 0.070 41.510 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 41.720 0.070 41.790 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 48.160 0.070 48.230 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 48.440 0.070 48.510 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 48.720 0.070 48.790 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 49.000 0.070 49.070 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 49.280 0.070 49.350 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 49.560 0.070 49.630 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 56.000 0.070 56.070 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 56.280 0.070 56.350 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal18 ;
      RECT 0.000 56.560 0.070 56.630 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal17 ;
      RECT 2.660 2.800 2.940 58.800 ;
      RECT 7.140 2.800 7.420 58.800 ;
      RECT 11.620 2.800 11.900 58.800 ;
      RECT 16.100 2.800 16.380 58.800 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal17 ;
      RECT 4.900 2.800 5.180 58.800 ;
      RECT 9.380 2.800 9.660 58.800 ;
      RECT 13.860 2.800 14.140 58.800 ;
    END
  END VDD
  OBS
    LAYER metal20 ;
    RECT 0 0 20.140 61.600 ;
    LAYER metal19 ;
    RECT 0 0 20.140 61.600 ;
    LAYER metal18 ;
    RECT 0.070 0 20.140 61.600 ;
    RECT 0 0.000 0.070 2.800 ;
    RECT 0 2.870 0.070 3.080 ;
    RECT 0 3.150 0.070 3.360 ;
    RECT 0 3.430 0.070 3.640 ;
    RECT 0 3.710 0.070 3.920 ;
    RECT 0 3.990 0.070 4.200 ;
    RECT 0 4.270 0.070 4.480 ;
    RECT 0 4.550 0.070 4.760 ;
    RECT 0 4.830 0.070 5.040 ;
    RECT 0 5.110 0.070 5.320 ;
    RECT 0 5.390 0.070 5.600 ;
    RECT 0 5.670 0.070 5.880 ;
    RECT 0 5.950 0.070 6.160 ;
    RECT 0 6.230 0.070 6.440 ;
    RECT 0 6.510 0.070 6.720 ;
    RECT 0 6.790 0.070 7.000 ;
    RECT 0 7.070 0.070 7.280 ;
    RECT 0 7.350 0.070 7.560 ;
    RECT 0 7.630 0.070 7.840 ;
    RECT 0 7.910 0.070 8.120 ;
    RECT 0 8.190 0.070 8.400 ;
    RECT 0 8.470 0.070 8.680 ;
    RECT 0 8.750 0.070 8.960 ;
    RECT 0 9.030 0.070 9.240 ;
    RECT 0 9.310 0.070 9.520 ;
    RECT 0 9.590 0.070 9.800 ;
    RECT 0 9.870 0.070 10.080 ;
    RECT 0 10.150 0.070 10.360 ;
    RECT 0 10.430 0.070 10.640 ;
    RECT 0 10.710 0.070 10.920 ;
    RECT 0 10.990 0.070 11.200 ;
    RECT 0 11.270 0.070 11.480 ;
    RECT 0 11.550 0.070 17.920 ;
    RECT 0 17.990 0.070 18.200 ;
    RECT 0 18.270 0.070 18.480 ;
    RECT 0 18.550 0.070 18.760 ;
    RECT 0 18.830 0.070 19.040 ;
    RECT 0 19.110 0.070 19.320 ;
    RECT 0 19.390 0.070 19.600 ;
    RECT 0 19.670 0.070 19.880 ;
    RECT 0 19.950 0.070 20.160 ;
    RECT 0 20.230 0.070 20.440 ;
    RECT 0 20.510 0.070 20.720 ;
    RECT 0 20.790 0.070 21.000 ;
    RECT 0 21.070 0.070 21.280 ;
    RECT 0 21.350 0.070 21.560 ;
    RECT 0 21.630 0.070 21.840 ;
    RECT 0 21.910 0.070 22.120 ;
    RECT 0 22.190 0.070 22.400 ;
    RECT 0 22.470 0.070 22.680 ;
    RECT 0 22.750 0.070 22.960 ;
    RECT 0 23.030 0.070 23.240 ;
    RECT 0 23.310 0.070 23.520 ;
    RECT 0 23.590 0.070 23.800 ;
    RECT 0 23.870 0.070 24.080 ;
    RECT 0 24.150 0.070 24.360 ;
    RECT 0 24.430 0.070 24.640 ;
    RECT 0 24.710 0.070 24.920 ;
    RECT 0 24.990 0.070 25.200 ;
    RECT 0 25.270 0.070 25.480 ;
    RECT 0 25.550 0.070 25.760 ;
    RECT 0 25.830 0.070 26.040 ;
    RECT 0 26.110 0.070 26.320 ;
    RECT 0 26.390 0.070 26.600 ;
    RECT 0 26.670 0.070 33.040 ;
    RECT 0 33.110 0.070 33.320 ;
    RECT 0 33.390 0.070 33.600 ;
    RECT 0 33.670 0.070 33.880 ;
    RECT 0 33.950 0.070 34.160 ;
    RECT 0 34.230 0.070 34.440 ;
    RECT 0 34.510 0.070 34.720 ;
    RECT 0 34.790 0.070 35.000 ;
    RECT 0 35.070 0.070 35.280 ;
    RECT 0 35.350 0.070 35.560 ;
    RECT 0 35.630 0.070 35.840 ;
    RECT 0 35.910 0.070 36.120 ;
    RECT 0 36.190 0.070 36.400 ;
    RECT 0 36.470 0.070 36.680 ;
    RECT 0 36.750 0.070 36.960 ;
    RECT 0 37.030 0.070 37.240 ;
    RECT 0 37.310 0.070 37.520 ;
    RECT 0 37.590 0.070 37.800 ;
    RECT 0 37.870 0.070 38.080 ;
    RECT 0 38.150 0.070 38.360 ;
    RECT 0 38.430 0.070 38.640 ;
    RECT 0 38.710 0.070 38.920 ;
    RECT 0 38.990 0.070 39.200 ;
    RECT 0 39.270 0.070 39.480 ;
    RECT 0 39.550 0.070 39.760 ;
    RECT 0 39.830 0.070 40.040 ;
    RECT 0 40.110 0.070 40.320 ;
    RECT 0 40.390 0.070 40.600 ;
    RECT 0 40.670 0.070 40.880 ;
    RECT 0 40.950 0.070 41.160 ;
    RECT 0 41.230 0.070 41.440 ;
    RECT 0 41.510 0.070 41.720 ;
    RECT 0 41.790 0.070 48.160 ;
    RECT 0 48.230 0.070 48.440 ;
    RECT 0 48.510 0.070 48.720 ;
    RECT 0 48.790 0.070 49.000 ;
    RECT 0 49.070 0.070 49.280 ;
    RECT 0 49.350 0.070 49.560 ;
    RECT 0 49.630 0.070 56.000 ;
    RECT 0 56.070 0.070 56.280 ;
    RECT 0 56.350 0.070 56.560 ;
    RECT 0 56.630 0.070 61.600 ;
    LAYER metal17 ;
    RECT 0 0 20.140 2.800 ;
    RECT 0 58.800 20.140 61.600 ;
    RECT 0.000 2.800 2.660 58.800 ;
    RECT 2.940 2.800 4.900 58.800 ;
    RECT 5.180 2.800 7.140 58.800 ;
    RECT 7.420 2.800 9.380 58.800 ;
    RECT 9.660 2.800 11.620 58.800 ;
    RECT 11.900 2.800 13.860 58.800 ;
    RECT 14.140 2.800 16.100 58.800 ;
    RECT 16.380 2.800 20.140 58.800 ;
  END
END fakeram45_64x32_upper

END LIBRARY
